module bnot(
    input logic a,
    output logic r
);

    assign r = ~a;

endmodule