module ram256x8();

endmodule