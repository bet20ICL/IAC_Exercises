module goodbye_world();
    initial begin
        $display("Goodbye bro");
    end
endmodule