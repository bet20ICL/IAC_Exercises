module hello_world();

    initial begin
        $display("Hello World");
        $fatal;
    end

endmodule